module washing_counter(
    input wire clk,
    input wire rst_n,
    input wire soft_rst,
    input wire start_washing,
    input wire [1:0] clk_freq,
    input wire round2_washing,
    output wire Washing_done 
);
reg [31:0] stop_count;
localparam [31:0] temp = 3'b100;
always @ *
begin
    case(clk_freq)
        2'b00: stop_count ='h11E1A300; 
        2'b01: stop_count = 'h23C34600;
        2'b10: stop_count = 'h47868C00;
        2'b11: stop_count = 'hFA56EA00;
    endcase
end    
reg [31:0] q;
always @(posedge clk or negedge rst_n) 
begin
    if(~rst_n)
        q <= 0;
    else if (~soft_rst)
        q <= 0;  
    else if (start_washing && ~Washing_done)
        q <= q + 1;
    else if (round2_washing)
    q <= 1;            
end
assign Washing_done = (q == stop_count);
endmodule